module delay #(
    parameter int CYCLES = 4, 
    parameter int 
)