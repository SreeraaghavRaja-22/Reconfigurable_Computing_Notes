package alu_pkg;
    typedef enum logic [1:0]{
        ADD_SEL = 2'b00,
        SUB_SEL = 2'b01,
        AND_SEL = 2'b10, 
        OR_SEL  = 2'b11
    } alu_sel_t;
endpackage